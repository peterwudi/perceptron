// megafunction wizard: %ALTMULT_ADD%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTMULT_ADD 

// ============================================================
// File Name: multAdd.v
// Megafunction Name(s):
// 			ALTMULT_ADD
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.0.1 Build 232 06/12/2013 SP 1 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module multAdd (
	dataa_0,
	dataa_1,
	dataa_2,
	dataa_3,
	datab_0,
	datab_1,
	datab_2,
	datab_3,
	result);

	input	[2:0]  dataa_0;
	input	[2:0]  dataa_1;
	input	[2:0]  dataa_2;
	input	[2:0]  dataa_3;
	input	[1:0]  datab_0;
	input	[1:0]  datab_1;
	input	[1:0]  datab_2;
	input	[1:0]  datab_3;
	output	[5:0]  result;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri0	[2:0]  dataa_0;
	tri0	[2:0]  dataa_1;
	tri0	[2:0]  dataa_2;
	tri0	[2:0]  dataa_3;
	tri0	[1:0]  datab_0;
	tri0	[1:0]  datab_1;
	tri0	[1:0]  datab_2;
	tri0	[1:0]  datab_3;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire [5:0] sub_wire0;
	wire [1:0] sub_wire10 = datab_3[1:0];
	wire [1:0] sub_wire9 = datab_2[1:0];
	wire [1:0] sub_wire8 = datab_1[1:0];
	wire [2:0] sub_wire5 = dataa_3[2:0];
	wire [2:0] sub_wire4 = dataa_2[2:0];
	wire [2:0] sub_wire3 = dataa_1[2:0];
	wire [5:0] result = sub_wire0[5:0];
	wire [2:0] sub_wire1 = dataa_0[2:0];
	wire [11:0] sub_wire2 = {sub_wire5, sub_wire4, sub_wire3, sub_wire1};
	wire [1:0] sub_wire6 = datab_0[1:0];
	wire [7:0] sub_wire7 = {sub_wire10, sub_wire9, sub_wire8, sub_wire6};

	altmult_add	ALTMULT_ADD_component (
				.dataa (sub_wire2),
				.datab (sub_wire7),
				.result (sub_wire0),
				.accum_sload (1'b0),
				.aclr0 (1'b0),
				.aclr1 (1'b0),
				.aclr2 (1'b0),
				.aclr3 (1'b0),
				.addnsub1 (1'b1),
				.addnsub1_round (1'b0),
				.addnsub3 (1'b1),
				.addnsub3_round (1'b0),
				.chainin (1'b0),
				.chainout_round (1'b0),
				.chainout_sat_overflow (),
				.chainout_saturate (1'b0),
				.clock0 (1'b1),
				.clock1 (1'b1),
				.clock2 (1'b1),
				.clock3 (1'b1),
				.coefsel0 ({3{1'b0}}),
				.coefsel1 ({3{1'b0}}),
				.coefsel2 ({3{1'b0}}),
				.coefsel3 ({3{1'b0}}),
				.datac ({88{1'b0}}),
				.ena0 (1'b1),
				.ena1 (1'b1),
				.ena2 (1'b1),
				.ena3 (1'b1),
				.mult01_round (1'b0),
				.mult01_saturation (1'b0),
				.mult0_is_saturated (),
				.mult1_is_saturated (),
				.mult23_round (1'b0),
				.mult23_saturation (1'b0),
				.mult2_is_saturated (),
				.mult3_is_saturated (),
				.output_round (1'b0),
				.output_saturate (1'b0),
				.overflow (),
				.rotate (1'b0),
				.scanina ({3{1'b0}}),
				.scaninb ({2{1'b0}}),
				.scanouta (),
				.scanoutb (),
				.shift_right (1'b0),
				.signa (1'b0),
				.signb (1'b0),
				.sourcea ({4{1'b0}}),
				.sourceb ({4{1'b0}}),
				.zero_chainout (1'b0),
				.zero_loopback (1'b0));
	defparam
		ALTMULT_ADD_component.accumulator = "NO",
		ALTMULT_ADD_component.addnsub_multiplier_pipeline_register1 = "UNREGISTERED",
		ALTMULT_ADD_component.addnsub_multiplier_pipeline_register3 = "UNREGISTERED",
		ALTMULT_ADD_component.addnsub_multiplier_register1 = "UNREGISTERED",
		ALTMULT_ADD_component.addnsub_multiplier_register3 = "UNREGISTERED",
		ALTMULT_ADD_component.chainout_adder = "NO",
		ALTMULT_ADD_component.chainout_register = "UNREGISTERED",
		ALTMULT_ADD_component.dedicated_multiplier_circuitry = "YES",
		ALTMULT_ADD_component.input_register_a0 = "UNREGISTERED",
		ALTMULT_ADD_component.input_register_a1 = "UNREGISTERED",
		ALTMULT_ADD_component.input_register_a2 = "UNREGISTERED",
		ALTMULT_ADD_component.input_register_a3 = "UNREGISTERED",
		ALTMULT_ADD_component.input_register_b0 = "UNREGISTERED",
		ALTMULT_ADD_component.input_register_b1 = "UNREGISTERED",
		ALTMULT_ADD_component.input_register_b2 = "UNREGISTERED",
		ALTMULT_ADD_component.input_register_b3 = "UNREGISTERED",
		ALTMULT_ADD_component.input_source_a0 = "DATAA",
		ALTMULT_ADD_component.input_source_a1 = "DATAA",
		ALTMULT_ADD_component.input_source_a2 = "DATAA",
		ALTMULT_ADD_component.input_source_a3 = "DATAA",
		ALTMULT_ADD_component.input_source_b0 = "DATAB",
		ALTMULT_ADD_component.input_source_b1 = "DATAB",
		ALTMULT_ADD_component.input_source_b2 = "DATAB",
		ALTMULT_ADD_component.input_source_b3 = "DATAB",
		ALTMULT_ADD_component.intended_device_family = "Stratix IV",
		ALTMULT_ADD_component.lpm_type = "altmult_add",
		ALTMULT_ADD_component.multiplier1_direction = "ADD",
		ALTMULT_ADD_component.multiplier3_direction = "ADD",
		ALTMULT_ADD_component.multiplier_register0 = "UNREGISTERED",
		ALTMULT_ADD_component.multiplier_register1 = "UNREGISTERED",
		ALTMULT_ADD_component.multiplier_register2 = "UNREGISTERED",
		ALTMULT_ADD_component.multiplier_register3 = "UNREGISTERED",
		ALTMULT_ADD_component.number_of_multipliers = 4,
		ALTMULT_ADD_component.output_register = "UNREGISTERED",
		ALTMULT_ADD_component.port_addnsub1 = "PORT_UNUSED",
		ALTMULT_ADD_component.port_addnsub3 = "PORT_UNUSED",
		ALTMULT_ADD_component.port_signa = "PORT_UNUSED",
		ALTMULT_ADD_component.port_signb = "PORT_UNUSED",
		ALTMULT_ADD_component.representation_a = "SIGNED",
		ALTMULT_ADD_component.representation_b = "SIGNED",
		ALTMULT_ADD_component.signed_pipeline_register_a = "UNREGISTERED",
		ALTMULT_ADD_component.signed_pipeline_register_b = "UNREGISTERED",
		ALTMULT_ADD_component.signed_register_a = "UNREGISTERED",
		ALTMULT_ADD_component.signed_register_b = "UNREGISTERED",
		ALTMULT_ADD_component.width_a = 3,
		ALTMULT_ADD_component.width_b = 2,
		ALTMULT_ADD_component.width_chainin = 1,
		ALTMULT_ADD_component.width_result = 6,
		ALTMULT_ADD_component.zero_chainout_output_register = "UNREGISTERED",
		ALTMULT_ADD_component.zero_loopback_output_register = "UNREGISTERED",
		ALTMULT_ADD_component.zero_loopback_pipeline_register = "UNREGISTERED",
		ALTMULT_ADD_component.zero_loopback_register = "UNREGISTERED";


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ACCUM_DIRECTION STRING "Add"
// Retrieval info: PRIVATE: ACCUM_SLOAD_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPE_REG STRING "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_REG STRING "0"
// Retrieval info: PRIVATE: ADDNSUB1_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ADDNSUB1_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB1_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ADDNSUB1_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB1_PIPE_REG STRING "0"
// Retrieval info: PRIVATE: ADDNSUB1_REG STRING "0"
// Retrieval info: PRIVATE: ADDNSUB3_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ADDNSUB3_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB3_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ADDNSUB3_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB3_PIPE_REG STRING "0"
// Retrieval info: PRIVATE: ADDNSUB3_REG STRING "0"
// Retrieval info: PRIVATE: ADD_ENABLE NUMERIC "0"
// Retrieval info: PRIVATE: ALL_REG_ACLR NUMERIC "0"
// Retrieval info: PRIVATE: A_ACLR_SRC_MULT0 NUMERIC "3"
// Retrieval info: PRIVATE: A_CLK_SRC_MULT0 NUMERIC "0"
// Retrieval info: PRIVATE: B_ACLR_SRC_MULT0 NUMERIC "3"
// Retrieval info: PRIVATE: B_CLK_SRC_MULT0 NUMERIC "0"
// Retrieval info: PRIVATE: CHAINOUT_OUTPUT_ACLR NUMERIC "3"
// Retrieval info: PRIVATE: CHAINOUT_OUTPUT_REG STRING "0"
// Retrieval info: PRIVATE: CHAINOUT_OUTPUT_REGISTER NUMERIC "0"
// Retrieval info: PRIVATE: CHAINOUT_OUTPUT_REGISTERED NUMERIC "0"
// Retrieval info: PRIVATE: CHAS_ZERO_CHAINOUT NUMERIC "0"
// Retrieval info: PRIVATE: HAS_ACCUMULATOR NUMERIC "0"
// Retrieval info: PRIVATE: HAS_ACUMM_SLOAD NUMERIC "0"
// Retrieval info: PRIVATE: HAS_CHAININ_PORT NUMERIC "0"
// Retrieval info: PRIVATE: HAS_CHAINOUT_ADDER NUMERIC "0"
// Retrieval info: PRIVATE: HAS_LOOPBACK NUMERIC "0"
// Retrieval info: PRIVATE: HAS_MAC STRING "0"
// Retrieval info: PRIVATE: HAS_SAT_ROUND STRING "0"
// Retrieval info: PRIVATE: HAS_ZERO_LOOPBACK NUMERIC "0"
// Retrieval info: PRIVATE: IMPL_STYLE_DEDICATED NUMERIC "1"
// Retrieval info: PRIVATE: IMPL_STYLE_DEFAULT NUMERIC "0"
// Retrieval info: PRIVATE: IMPL_STYLE_LCELL NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
// Retrieval info: PRIVATE: MULT_REGA0 NUMERIC "0"
// Retrieval info: PRIVATE: MULT_REGB0 NUMERIC "0"
// Retrieval info: PRIVATE: MULT_REGOUT0 NUMERIC "0"
// Retrieval info: PRIVATE: NUM_MULT STRING "4"
// Retrieval info: PRIVATE: OP1 STRING "Add"
// Retrieval info: PRIVATE: OP3 STRING "Add"
// Retrieval info: PRIVATE: OUTPUT_EXTRA_LAT NUMERIC "0"
// Retrieval info: PRIVATE: OUTPUT_REG_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: OUTPUT_REG_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: Q_ACLR_SRC_MULT0 NUMERIC "3"
// Retrieval info: PRIVATE: Q_CLK_SRC_MULT0 NUMERIC "0"
// Retrieval info: PRIVATE: REG_OUT NUMERIC "0"
// Retrieval info: PRIVATE: RNFORMAT STRING "6"
// Retrieval info: PRIVATE: ROTATE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROTATE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROTATE_OUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROTATE_OUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROTATE_OUT_REG STRING "0"
// Retrieval info: PRIVATE: ROTATE_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROTATE_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROTATE_PIPE_REG STRING "0"
// Retrieval info: PRIVATE: ROTATE_REG STRING "0"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_MODE STRING "Enabled"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_OUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_OUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_OUT_REG STRING "0"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_PIPE_REG STRING "0"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_REG STRING "0"
// Retrieval info: PRIVATE: ROUND3_FRAC_WIDTH NUMERIC "-1"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_CHAINOUT_TYPE STRING "Nearest Integer"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_MODE STRING "Disabled"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_PIPE_REG STRING "0"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_REG STRING "0"
// Retrieval info: PRIVATE: RQFORMAT STRING "Q1.15"
// Retrieval info: PRIVATE: RTS_WIDTH STRING "6"
// Retrieval info: PRIVATE: SAME_CONFIG NUMERIC "1"
// Retrieval info: PRIVATE: SAME_CONTROL_SRC_A0 NUMERIC "1"
// Retrieval info: PRIVATE: SAME_CONTROL_SRC_B0 NUMERIC "1"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_MODE STRING "Enabled"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_OUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_OUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_PIPE_REG STRING "0"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_REG STRING "0"
// Retrieval info: PRIVATE: SAT3_FRAC_WIDTH NUMERIC "2"
// Retrieval info: PRIVATE: SAT3_OUTPUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SAT3_OUTPUT_CHAINOUT_TYPE STRING "Asymmetric"
// Retrieval info: PRIVATE: SAT3_OUTPUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_OUTPUT_MODE STRING "Enabled"
// Retrieval info: PRIVATE: SAT3_OUTPUT_OVERFLOW NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_OUTPUT_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SAT3_OUTPUT_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_OUTPUT_PIPE_REG STRING "0"
// Retrieval info: PRIVATE: SAT3_OUTPUT_REG STRING "0"
// Retrieval info: PRIVATE: SCANOUTA NUMERIC "0"
// Retrieval info: PRIVATE: SCANOUTB NUMERIC "0"
// Retrieval info: PRIVATE: SHIFTOUTA_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SHIFTOUTA_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SHIFTOUTA_REG STRING "0"
// Retrieval info: PRIVATE: SHIFT_RIGHT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SHIFT_RIGHT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SHIFT_RIGHT_OUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SHIFT_RIGHT_OUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SHIFT_RIGHT_OUT_REG STRING "0"
// Retrieval info: PRIVATE: SHIFT_RIGHT_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SHIFT_RIGHT_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SHIFT_RIGHT_PIPE_REG STRING "0"
// Retrieval info: PRIVATE: SHIFT_RIGHT_REG STRING "0"
// Retrieval info: PRIVATE: SHIFT_ROTATE_MODE STRING "None"
// Retrieval info: PRIVATE: SIGNA STRING "SIGNED"
// Retrieval info: PRIVATE: SIGNA_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SIGNA_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SIGNA_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SIGNA_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SIGNA_PIPE_REG STRING "0"
// Retrieval info: PRIVATE: SIGNA_REG STRING "0"
// Retrieval info: PRIVATE: SIGNB STRING "SIGNED"
// Retrieval info: PRIVATE: SIGNB_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SIGNB_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SIGNB_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SIGNB_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SIGNB_PIPE_REG STRING "0"
// Retrieval info: PRIVATE: SIGNB_REG STRING "0"
// Retrieval info: PRIVATE: SRCA0 STRING "Multiplier input"
// Retrieval info: PRIVATE: SRCB0 STRING "Multiplier input"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: WIDTHA STRING "3"
// Retrieval info: PRIVATE: WIDTHB STRING "2"
// Retrieval info: PRIVATE: ZERO_CHAINOUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ZERO_CHAINOUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ZERO_CHAINOUT_REG STRING "0"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_OUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_OUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_OUT_REG STRING "0"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_PIPE_REG STRING "0"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_REG STRING "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: ACCUMULATOR STRING "NO"
// Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_PIPELINE_REGISTER1 STRING "UNREGISTERED"
// Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_PIPELINE_REGISTER3 STRING "UNREGISTERED"
// Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_REGISTER1 STRING "UNREGISTERED"
// Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_REGISTER3 STRING "UNREGISTERED"
// Retrieval info: CONSTANT: CHAINOUT_ADDER STRING "NO"
// Retrieval info: CONSTANT: CHAINOUT_REGISTER STRING "UNREGISTERED"
// Retrieval info: CONSTANT: DEDICATED_MULTIPLIER_CIRCUITRY STRING "YES"
// Retrieval info: CONSTANT: INPUT_REGISTER_A0 STRING "UNREGISTERED"
// Retrieval info: CONSTANT: INPUT_REGISTER_A1 STRING "UNREGISTERED"
// Retrieval info: CONSTANT: INPUT_REGISTER_A2 STRING "UNREGISTERED"
// Retrieval info: CONSTANT: INPUT_REGISTER_A3 STRING "UNREGISTERED"
// Retrieval info: CONSTANT: INPUT_REGISTER_B0 STRING "UNREGISTERED"
// Retrieval info: CONSTANT: INPUT_REGISTER_B1 STRING "UNREGISTERED"
// Retrieval info: CONSTANT: INPUT_REGISTER_B2 STRING "UNREGISTERED"
// Retrieval info: CONSTANT: INPUT_REGISTER_B3 STRING "UNREGISTERED"
// Retrieval info: CONSTANT: INPUT_SOURCE_A0 STRING "DATAA"
// Retrieval info: CONSTANT: INPUT_SOURCE_A1 STRING "DATAA"
// Retrieval info: CONSTANT: INPUT_SOURCE_A2 STRING "DATAA"
// Retrieval info: CONSTANT: INPUT_SOURCE_A3 STRING "DATAA"
// Retrieval info: CONSTANT: INPUT_SOURCE_B0 STRING "DATAB"
// Retrieval info: CONSTANT: INPUT_SOURCE_B1 STRING "DATAB"
// Retrieval info: CONSTANT: INPUT_SOURCE_B2 STRING "DATAB"
// Retrieval info: CONSTANT: INPUT_SOURCE_B3 STRING "DATAB"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altmult_add"
// Retrieval info: CONSTANT: MULTIPLIER1_DIRECTION STRING "ADD"
// Retrieval info: CONSTANT: MULTIPLIER3_DIRECTION STRING "ADD"
// Retrieval info: CONSTANT: MULTIPLIER_REGISTER0 STRING "UNREGISTERED"
// Retrieval info: CONSTANT: MULTIPLIER_REGISTER1 STRING "UNREGISTERED"
// Retrieval info: CONSTANT: MULTIPLIER_REGISTER2 STRING "UNREGISTERED"
// Retrieval info: CONSTANT: MULTIPLIER_REGISTER3 STRING "UNREGISTERED"
// Retrieval info: CONSTANT: NUMBER_OF_MULTIPLIERS NUMERIC "4"
// Retrieval info: CONSTANT: OUTPUT_REGISTER STRING "UNREGISTERED"
// Retrieval info: CONSTANT: PORT_ADDNSUB1 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_ADDNSUB3 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_SIGNA STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_SIGNB STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: REPRESENTATION_A STRING "SIGNED"
// Retrieval info: CONSTANT: REPRESENTATION_B STRING "SIGNED"
// Retrieval info: CONSTANT: SIGNED_PIPELINE_REGISTER_A STRING "UNREGISTERED"
// Retrieval info: CONSTANT: SIGNED_PIPELINE_REGISTER_B STRING "UNREGISTERED"
// Retrieval info: CONSTANT: SIGNED_REGISTER_A STRING "UNREGISTERED"
// Retrieval info: CONSTANT: SIGNED_REGISTER_B STRING "UNREGISTERED"
// Retrieval info: CONSTANT: WIDTH_A NUMERIC "3"
// Retrieval info: CONSTANT: WIDTH_B NUMERIC "2"
// Retrieval info: CONSTANT: WIDTH_CHAININ NUMERIC "1"
// Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "6"
// Retrieval info: CONSTANT: ZERO_CHAINOUT_OUTPUT_REGISTER STRING "UNREGISTERED"
// Retrieval info: CONSTANT: ZERO_LOOPBACK_OUTPUT_REGISTER STRING "UNREGISTERED"
// Retrieval info: CONSTANT: ZERO_LOOPBACK_PIPELINE_REGISTER STRING "UNREGISTERED"
// Retrieval info: CONSTANT: ZERO_LOOPBACK_REGISTER STRING "UNREGISTERED"
// Retrieval info: USED_PORT: dataa_0 0 0 3 0 INPUT GND "dataa_0[2..0]"
// Retrieval info: USED_PORT: dataa_1 0 0 3 0 INPUT GND "dataa_1[2..0]"
// Retrieval info: USED_PORT: dataa_2 0 0 3 0 INPUT GND "dataa_2[2..0]"
// Retrieval info: USED_PORT: dataa_3 0 0 3 0 INPUT GND "dataa_3[2..0]"
// Retrieval info: USED_PORT: datab_0 0 0 2 0 INPUT GND "datab_0[1..0]"
// Retrieval info: USED_PORT: datab_1 0 0 2 0 INPUT GND "datab_1[1..0]"
// Retrieval info: USED_PORT: datab_2 0 0 2 0 INPUT GND "datab_2[1..0]"
// Retrieval info: USED_PORT: datab_3 0 0 2 0 INPUT GND "datab_3[1..0]"
// Retrieval info: USED_PORT: result 0 0 6 0 OUTPUT GND "result[5..0]"
// Retrieval info: CONNECT: @dataa 0 0 3 0 dataa_0 0 0 3 0
// Retrieval info: CONNECT: @dataa 0 0 3 3 dataa_1 0 0 3 0
// Retrieval info: CONNECT: @dataa 0 0 3 6 dataa_2 0 0 3 0
// Retrieval info: CONNECT: @dataa 0 0 3 9 dataa_3 0 0 3 0
// Retrieval info: CONNECT: @datab 0 0 2 0 datab_0 0 0 2 0
// Retrieval info: CONNECT: @datab 0 0 2 2 datab_1 0 0 2 0
// Retrieval info: CONNECT: @datab 0 0 2 4 datab_2 0 0 2 0
// Retrieval info: CONNECT: @datab 0 0 2 6 datab_3 0 0 2 0
// Retrieval info: CONNECT: result 0 0 6 0 @result 0 0 6 0
// Retrieval info: GEN_FILE: TYPE_NORMAL multAdd.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL multAdd.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL multAdd.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL multAdd.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL multAdd_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL multAdd_bb.v FALSE
// Retrieval info: LIB_FILE: altera_mf
